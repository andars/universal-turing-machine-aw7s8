`default_nettype none

module user_module_341174563322724948(
  input [7:0] io_in,
  output [7:0] io_out
);

// TODO
assign io_out[0] = ~io_in[0];
assign io_out[1] = ~io_in[0];

endmodule
